class transaction;
  rand bit in1;
  bit out;
  constraint in_c{in1 inside {[0:1]};}
endclass

  
