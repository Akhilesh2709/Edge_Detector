interface add_if(input logic clk,reset);
  logic in1;
  logic out;
endinterface
